// Author: Colin Pollard, Ian Lavin
// Date: 10/15/2020
// This file creates an FSM to control basic R-type instructions.

module R_Type_FSM(clk, rst, dataInA, dataInB, addressA, addressB, weA, weB, dataOutA, dataOutB);
input clk;



endmodule