/*
 * Author: Colin Pollard, Ian Lavin, Luke Majors, Mckay Mower
 * Date: 9/17/2020
 *
 * This module represents a finite state machine that is used to test the ALU
 * and the register file. This fsm specifically computes a fibonacci sequence
 * using the ALU and regfile.
 */
 
 //module fib_test_fsm(clk, rst, reg_write, regA, regB, op, reg_imm, 